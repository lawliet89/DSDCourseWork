fp_add_sub_inst : fp_add_sub PORT MAP (
		add_sub	 => add_sub_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
