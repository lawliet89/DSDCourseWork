const_7_inst : const_7 PORT MAP (
		result	 => result_sig
	);
